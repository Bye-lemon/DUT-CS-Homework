library verilog;
use verilog.vl_types.all;
entity FIFO_vlg_vec_tst is
end FIFO_vlg_vec_tst;
