LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CNT4 IS                              -- 8λ���Լ��ؼӷ�������
    PORT (    CLK 		: IN STD_LOGIC;
					Q	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END CNT4;
ARCHITECTURE behav OF CNT4 IS
    SIGNAL COUNT : STD_LOGIC_VECTOR (3 DOWNTO 0);
BEGIN
    PROCESS( CLK )
    BEGIN
        IF CLK'EVENT AND CLK = '1' THEN
           COUNT <= COUNT + 1;
        END IF;
		Q  <= COUNT;
    END PROCESS;
END behav;

