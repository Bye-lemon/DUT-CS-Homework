library verilog;
use verilog.vl_types.all;
entity CNT10_vlg_vec_tst is
end CNT10_vlg_vec_tst;
