library verilog;
use verilog.vl_types.all;
entity ROM_vlg_vec_tst is
end ROM_vlg_vec_tst;
